module multiplier ( 
    
    // Inputs
    input wire clk_i,
    input wire rst_i,
    input wire [31:0] op_A_i,
    input wire [31:0] op_B_i,
    input wire ext_A_i,
    input wire ext_B_i,
    input wire upper_i,

    // Outputs
    output wire [31:0] result_o,
    output done_o
);

// CONTROL PATH

// DATA PATH

endmodule